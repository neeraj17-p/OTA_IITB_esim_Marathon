.title KiCad schematic
U1 OUT plot_v1
M4 OUT M34G VDD VDD pmos
M2 OUT VINN ID5 GND nmos
M1 M34G VINP ID5 GND nmos
VDD1 VDD GND DC 
M3 M34G M34G VDD VDD pmos
Vbias1 VBIAS GND DC 
VINP1 VINP GND DC 
VINN1 VINN GND DC 
M5 ID5 VBIAS GND GND nmos
.end
