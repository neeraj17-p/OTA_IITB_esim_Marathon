.title KiCad schematic
vinp1 VINP NODEP AC
M6 SOURCETAIL VBCAS MSD GND nmos
vbcas1 VBCAS GND DC
M1 DRAINL VINP SOURCETAIL GND nmos
vinpb1 NODEP GND DC
M3 DRAINL DRAINL VDD VDD pmos
vdd1 VDD GND DC
M5 MSD VBIAS GND GND nmos
Itail1 GND SOURCETAIL dc
U1 OUT plot_db
CL1 OUT GND 5p
M4 OUT DRAINL VDD VDD pmos
M2 OUT VINN SOURCETAIL GND nmos
vinn1 VINN NODEN AC
vinnb1 NODEN GND DC
vbias1 VBIAS GND DC
.end
